package apb_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "afvip_apb_sequence_item.svh"
    `include "afvip_apb_sequencer.svh"
    `include "afvip_apb_driver.svh"
    `include "afvip_apb_monitor.svh"
    `include "afvip_apb_agent.svh"
    `include "afvip_apb_sequence.svh"
endpackage