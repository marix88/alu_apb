package rst_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "afvip_reset_sequence_item.svh"
    `include "afvip_reset_sequencer.svh"
    `include "afvip_reset_driver.svh"
    `include "afvip_reset_monitor.svh"
    `include "afvip_reset_agent.svh"
    `include "afvip_reset_sequence.svh"
endpackage