package intr_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "afvip_interrupt_sequence_item.svh"
    `include "afvip_interrupt_monitor.svh"
    `include "afvip_interrupt_agent.svh"  
endpackage