package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import apb_pkg::*;
    import intr_pkg::*;
    import rst_pkg::*;
    import env_scb_pkg::*;
    `include "afvip_test.svh"
endpackage