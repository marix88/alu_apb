package env_scb_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import apb_pkg::*;
    import intr_pkg::*;
    import rst_pkg::*;
    `include "afvip_scoreboard.svh" 
    `include "afvip_environment.svh" 
    //`include "afvip_coverage.svh"
endpackage